library verilog;
use verilog.vl_types.all;
entity CPUp1_vlg_vec_tst is
end CPUp1_vlg_vec_tst;
