library verilog;
use verilog.vl_types.all;
entity CPUp2_vlg_vec_tst is
end CPUp2_vlg_vec_tst;
