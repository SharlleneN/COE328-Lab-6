LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

entity ALU is -- ALU unit includes Reg. 3
port ( clk, reset : in std_logic ;
sign : out std_logic;
studentID : in std_logic_vector(3 downto 0); -- student number
Reg1, Reg2: in std_logic_vector(7 downto 0); -- 8-bit inputs A & B from Reg. 1 & Reg. 2
opcode : in std_logic_vector(7 downto 0); -- 8-bit opcode from Decoder
R1,R2,R3: out std_logic_vector(3 downto 0)); -- 4-bit Results
end ALU ;

architecture calculation of ALU is
SIGNAL result : STD_logic_Vector(9 downto 0);
SIGNAL temp1,temp2: STD_logic_Vector(3 downto 0);
begin
	process ( clk, reset )
		begin
			if reset = '1' then
			result <= "0000000000" ;
			elsif (clk'EVENT AND clk = '1') then
			case opcode is
					when "00000001" =>
					sign <= '0';
					result <= "00" & (Reg1 + Reg2);
					when "00000010" =>
					IF (Reg1(7 downto 0) >= Reg2(7 downto 0))THEN
					sign <= '0';
					result <= "00" & (Reg1 - Reg2);
					ELSE
					sign <= '1';
					result <= "00" & (Reg2 - Reg1);
					END IF;
					when "00000100" =>
					sign <= '0';
					result <= "00" & not(Reg1);
					when "00001000" =>
					sign <= '0';
					result <= "00" & not(Reg1 AND Reg2);
					when "00010000" =>
					sign <= '0';
					result <= "00" & not(Reg1 OR Reg2);
					when "00100000" =>
					sign <= '0';
					result <= "00" &(Reg1 AND Reg2);
					when "01000000" =>
					result <= "00" & (Reg1 XOR Reg2);
					when "10000000" =>
					sign <= '0';
					result <= "00" & (Reg1 OR Reg2);
					when others =>
					result <= "0000000000";
end case;
end if ;
end process ;

R1 <= result(3 downto 0);
R2 <= result(7 downto 4);
R3 <= studentID(3 downto 0);

end calculation;